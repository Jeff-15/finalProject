Blue
0 0 0 0 0 h 1 B 9 B 
0 0 0 0 0 h 3 B 11 B 
0 0 0 0 0 h 5 B 19 B 
0 0 0 0 0 h 7 B 21 B 
1 5 5 7 4 3 4 4 3 5 1 9 4 10 0 4 0 8 2 9 1 10 1 6 0 11 3 12 2 11 3 3 0 8 2 2 2 6 
14
