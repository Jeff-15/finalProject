Blue
0 0 0 0 0 h 1 B 13 B 
0 0 0 0 0 h 3 B 21 B 
0 0 0 0 0 h 5 B 25 B 
0 0 0 0 0 h 11 B 33 B 
